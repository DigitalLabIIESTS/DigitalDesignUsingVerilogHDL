`timescale 1ns / 1ps
module half_adder_struct(sum_out,carry_out,a_in,b_in);
    output sum_out;
    output carry_out;
    input a_in,b_in;
endmodule
